//或门逻辑描述
module or2a(a,b,c);
	input a,b;
	output c;
	assign c = a | b;
endmodule 