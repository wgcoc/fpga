//含义异步复位/时钟使能型触发器
//含异步清零和时钟同步使能得D触发起
module DFF2(CLK,D,Q,RST,EN);
	input CLK,D,RST,EN;
	output Q;
	reg Q;
	/*1.敏感信号表一旦含有posedge或negedge的边沿敏感信号后，
	    所有其它电平型敏感变量都不能放在敏感信号列表，从而导致此过程中所有这些
	    未能进入敏感信号表的变量都必须是相对于时钟同步
	  2.如果希望在同一模块中含有独立于主时钟的时序或逻辑，则必须用另一个过程来描述
	  3.如果某信号A被定义为边沿敏感时钟信号，则必须在敏感信号表中给出对应的表述，
	    如posedge A或negedge A；但在always过程结构中不能再出现信号A了
	  4.如果将某信号B定义为对应于时钟的电平敏感的异步控制信号（或仅仅是异步输入信号），
	    则除了在敏感信号表中给出对应的描述外，如posedge B或negedge B，在always过程
		 结构中必须明示信号B的逻辑行为，如本例的RST。特表注意这种表述的不一致性，即表述
		 上必须是边沿敏感信号，如posedge B，但电路性能上是电平敏感的
	  5.如果将某信号定义为对应于时钟的同步控制信号（或仅仅是同步输入信号），则绝不可以
	    以任何形式出现在敏感信号表中
	  6.敏感信号表中一旦出现类似posedge或negedge的边沿敏感信号，则不允许再出现其它
	    非敏感信号的报表述。即敏感和非敏感表述不能同时出现在敏感信号表中，每一个过程
		 语句只能放置一种类型的敏感信号，不能混放
	*/
	always @(posedge CLK,negedge RST)
	begin
		if(!RST) Q <= 0;		//如果RST=0条件成立，Q被清零
		else if(EN) Q <= D;	//在CLK上升沿处，EN=1，则执行赋值语句
 	end 
endmodule 