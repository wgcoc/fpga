//异步时序模块
/*1.在时序电路设计中应注意：一个时钟过程只能构成对应单一时钟信号的时序电路，
    如果在某一过程中需要构成多触发器时序电路，也只能产生对应某个单一时钟的同步时序逻辑
  2.没有单一主控时钟的时序电路（或系统）中所有的时序部件不随某个主控时钟同步接受时钟信号
    达到状态同步变化的电路都属于异步时序电路
  3.现代数字系统中，很少有应用异步时序逻辑的场合
*/
module AMOD(D,A,CLK,Q); //含有两个过程语句的异步时序电路
 	input A,D,CLK;
	output Q;
	reg Q,Q1;
	//过程1
	always @(posedge CLK)
	begin 
		Q1 = ~(A | Q);
	end
	//过程2，将过程1的输出作为时钟信号
	always @(posedge Q1)
	begin
		Q = D;
	end
endmodule 