module MUX41a_v3(A,B,C,D,S1,S0,Y);
	input A,B,C,D,S1,S0;
	output Y;
	//定义一个always@模块内部的暂存变量SEL[1:0]
	reg [1:0] SEL;
	//定义一个always@模块内部的输出端口信号
	reg Y;
	always @(A,B,C,D,SEL)
	begin //语句块起始
		SEL = {S1,S0}; //把S1,S0并位为2元素矢量变量SEL[1:0]
		/* 1.“=”表示阻塞赋值符号；“<=”表示非阻塞式赋值
			2.阻塞赋值的特点：如果在一个语句块中含有多条阻塞式赋值语句，
			  而当执行到其中某条赋值语句时，其他语句被禁止执行，这是其
			  他语句如同被阻塞了一样
			  非阻塞赋值的特点：必须在块语句执行结束时才整体完成赋值操作
			3.assign语句和always语句中出现的赋值符号“=”从理论上说是不同性质的，
			  因为前者属于连续赋值语句，具有并行赋值特性，后者属于过程赋值类中的
			  顺序赋值语句。但从综合角度看其结果是相同的。
		*/
		if(SEL == 0)		Y = A;
		else if(SEL == 1)	Y = B;
		else if(SEL == 2)	Y = C;
		else					Y = D;
	end
endmodule 